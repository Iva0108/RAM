`ifndef RAM_PKG
`define RAM_PKG

package ram_pkg;
	`include "transaction.sv"
	`include "generator.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "scoreboard.sv"
	`include "environment.sv"
endpackage

`endif